module instruction_mem(instruction, reset, im_readAddr);
	output [31:0] instruction;
	input [6:0] im_readAddr;
	input reset;
	
	reg [31:0] mem[127:0];
	
	assign mem[0] = 32'b00100000000100000000000000000111;
	assign mem[1] = 32'b00100000000010000000000000000111;
	assign mem[2] = 32'b10101110000010000000000000000000;
	assign mem[3] = 32'b10001110000010000000000000000000;
	
	assign mem[4] = 32'b00100000000100010000000000000101;
	assign mem[5] = 32'b00100000000010010000000000000101;
	assign mem[6] = 32'b10101110001010010000000000000000;
	assign mem[7] = 32'b10001110001010010000000000000000;
	
	assign mem[8] =  32'b00100000000100100000000000000011;
	assign mem[9] =  32'b00100000000010100000000000000011;
	assign mem[10] = 32'b10101110010010100000000000000000;
	assign mem[11] = 32'b10001110010010100000000000000000;
	 
	assign mem[12] = 32'b00100000000100110000000000000101;
	assign mem[13] = 32'b00100000000010110000000000000101;
	assign mem[14] = 32'b10101110011010110000000000000000;
	assign mem[15] = 32'b10001110011010110000000000000000;
	  
	assign mem[16] = 32'b00000010011000001100000000100000;
	  
	assign mem[17] = 32'b00100000000101000101101001011010;
	assign mem[18] = 32'b00100000000011000101101001011010;
	assign mem[19] = 32'b10101110100011000000000000000000;
	assign mem[20] = 32'b10001110100011000000000000000000;
	
	assign mem[21] = 32'b00100000000101010110011101100111;
	assign mem[22] = 32'b00100000000011010110011101100111;
	assign mem[23] = 32'b10101110101011010000000000000000;
	assign mem[24] = 32'b10001110101011010000000000000000;
	
	assign mem[25] = 32'b00100000000101100000000000111100;
	assign mem[26] = 32'b00100000000011100000000000111100;
	assign mem[27] = 32'b10101110110011100000000000000000;
	assign mem[28] = 32'b10001110110011100000000000000000;
	
	assign mem[29] = 32'b00100000000101110000000011111111;
	assign mem[30] = 32'b00100000000011110000000011111111;
	assign mem[31] = 32'b10101110111011110000000000000000;
	assign mem[32] = 32'b10001110111011110000000000000000;
	
	assign mem[33] = 32'b00000001000010010001000000100010;
	assign mem[34] = 32'b00100000000110010000000000000011;
	assign mem[35] = 32'b00011100010110010000000000000100;

	assign mem[36] = 32'b00000001010110010101000000000000;
	assign mem[37] = 32'b00100000000010110000000000000111;
	assign mem[38] = 32'b00000001100011010111000000100100;
	
	assign mem[39] = 32'b00001000000000000000000000101011;
	assign mem[40] = 32'b00100001010010100000000000000100;
	assign mem[41] = 32'b00000001010110010101100000100010;
	assign mem[42] = 32'b00000001100011010111000000100101;
	
	assign mem[43] = 32'b00000001000010010100000000100000;
	assign mem[44] = 32'b00000001100011010001100000100110;
	assign mem[45] = 32'b00000000011011110111000000100100;
	
	
	
	
	//assign instruction = reset ? mem[im_readAddr] : 32'b0;
	always@(*)
	if(reset)
	instruction <= mem[im_readAddr];
	else 
	instruction <= 32'b0;
endmodule
